import Vector::*;
import Randomizable::*;
import Multi::*;

(* synthesize *)
module mkTestReferenceMultiplier ();
endmodule 

(* synthesize *)
module mkTestSingleCycleMultiplier();
endmodule 
