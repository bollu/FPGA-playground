package FirstAttempt;
    module mkHelloWorld ();
        rule sayhello (True);
            $display("hello, world");
        endrule
    endmodule
endpackage
