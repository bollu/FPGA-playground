import Vector::*;
import Randomizable::*;
import Multi::*;

(* synthesize *)
module TestReferenceMultiplier 
endmodule 

(* synthesize *)
module TestSingleCycleMultiplier
endmodule 
